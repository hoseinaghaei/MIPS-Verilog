// `timescale 1ns / 1ps

////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer:
//
// Create Date:   13:20:00 07/21/2022
// Design Name:   FP_ALU
// Module Name:   E:/edu/term6/CA/phase4/Phase4/FP_ALU_test.v
// Project Name:  Phase4
// Target Device:  
// Tool versions:  
// Description: 
//
// Verilog Test Fixture created by ISE for module: FP_ALU
//
// Dependencies:
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
////////////////////////////////////////////////////////////////////////////////

module FP_ALU_test;

	// Inputs
	reg [31:0] num1;
	reg [31:0] num2;
	reg [2:0] func;

	// Outputs
	wire [31:0] result;
	wire overflow;
	wire underflow;
	wire inexact;
	wire div_by_zero;
	wire QNaN;
	wire SNaN;

	// Instantiate the Unit Under Test (UUT)
	FP_ALU uut (
		.num1(num1), 
		.num2(num2), 
		.func(func), 
		.result(result), 
		.overflow(overflow), 
		.underflow(underflow), 
		.inexact(inexact), 
		.div_by_zero(div_by_zero), 
		.QNaN(QNaN), 
		.SNaN(SNaN)
	);

	initial begin
		// Initialize Inputs
		num1 = 0;
		num2 = 0;
		func = 0;

		#10;    	
		// add test 
      num1 = 32'b01000001000001000000000000000000;
		num2 = 32'b00111111101000000000000000000000;
		func = 3'b000;
 //8.25+1.25=9.5 01000001000010000000000000000000
		
		#10;    	
		// add test 
      num1 = 32'b01000001000001000000000000000000;
		num2 = 32'b10111111101000000000000000000000;
		func = 3'b000;
 //8.25+-1.25=7  01000000111000000000000000000000
		 
		#10;    	
		// add test 
      num1 = 32'b11000001000001000000000000000000;
		num2 = 32'b10111111101000000000000000000000;
		func = 3'b000;
//-8.25+-1.25=-9.5 11000001000010000000000000000000
		
		#10;    	
		// add test 
      num1 = 32'b11000001000001000000000000000000;
		num2 = 32'b10111111101000000000000000000000;
		func = 3'b000;
//-8.25+1.25=-7 11000000111000000000000000000000

		#10;    	
		// add test 
      num1 = 32'b10111111101000000000000000000000;
		num2 = 32'b00111111101000000000000000000000;
		func = 3'b000;
 //-1.25+1.25=0  00000000000000000000000000000000	
		
		#10
		// add test inexact test
      num1 = 32'b01000001000001000000000000000000;
		num2 = 32'b10111111101000000000000000000001;
		func = 3'b000;
 //8.25+-1.25+eps=7  01000000111000000000000000000000
		
		#10;    	
		// add test 
      num1 = 32'b01111111100000000000000000000000;
		num2 = 32'b00111111101000000000000000000000;
		func = 3'b000;
 //inf+1.25=inf 01000001000010000000000000000000
 
		#10;    	
		// add test 
      num1 = 32'b11111111100000000000000000000000;
		num2 = 32'b00111111101000000000000000000000;
		func = 3'b000;
 //-inf+1.25=-inf 01000001000010000000000000000000
 
		#10;    	
		// add test 
      num1 = 32'b11111111100000000000000000000000;
		num2 = 32'b01111111100000000000000000000000;
		func = 3'b000;
 //-inf+inf=qnan 01000001000010000000000000000000
 
		#10;    	
		// sub test 
      num1 = 32'b01000001000001000000000000000000;
		num2 = 32'b00111111101000000000000000000000;
		func = 3'b001;
 //8.25-1.25=7 01000000111000000000000000000000 
		
		#10;    	
		// sub test 
      num1 = 32'b01000001000001000000000000000000;
		num2 = 32'b10111111101000000000000000000000;
		func = 3'b001;
 //8.25--1.25=9.5  01000001000010000000000000000000
		 
		#10;    	
		// sub test 
      num1 = 32'b11000001000001000000000000000000;
		num2 = 32'b10111111101000000000000000000000;
		func = 3'b001;
//-8.25--1.25=-7 11000000111000000000000000000000 
		
		#10;    	
		// sub test 
      num1 = 32'b11000001000001000000000000000000;
		num2 = 32'b10111111101000000000000000000000;
		func = 3'b001;
//-8.25-1.25=-9.5 11000001000010000000000000000000

		#10;    	
		// sub test 
      num1 = 32'b00111111101000000000000000000000;
		num2 = 32'b00111111101000000000000000000000;
		func = 3'b001;
 //1.25+1.25=0  00000000000000000000000000000000
		
		#10;    	
		// mul test 
      num1 = 32'b01000001000001000000000000000000;
		num2 = 32'b00111111101000000000000000000000;
		func = 3'b010;
 //8.25*1.25=10.3125  0_10000010_01001010000000000000000
		
		#10;
		// mul test 
      num1 = 32'b01000001000001000000000000000000;
		num2 = 32'b10111111101000000000000000000000;
		func = 3'b010;
 //8.25*-1.25=-10.3125  1_10000010_01001010000000000000000
		
		#10;
		// mul test 
      num1 = 32'b01000001000001000000000000000000;
		num2 = 32'b0;
		func = 3'b010;
 //8.25*0=0  0
		
		
		#10;    	
		// mul test 
      num1 = 32'b01111111100000000000000000000000;
		num2 = 32'b00111111101000000000000000000000;
		func = 3'b010;
 //inf*1.25=inf  0_10000010_01001010000000000000000
		
		#10; 
		// mul test 
      num1 = 32'b01111111100000000000000000000000;
		num2 = 32'b10111111101000000000000000000000;
		func = 3'b010;
 //inf*-1.25=-inf  0_10000010_01001010000000000000000
		
		#10; 
		// mul test 
      num1 = 32'b01111111100000000000000000000000;
		num2 = 32'b00000000000000000000000000000000;
		func = 3'b010;
 //inf*0=-qnan  0_10000010_01001010000000000000000
		
		
		#10;
		// div by zero test 
      num1 = 32'b01000001000001000000000000000000;
		num2 = 32'b0;
		func = 3'b011;
 //8.25/0=div by zero  0
		
		#10;
		// div test 
      num1 = 32'b01000001000001000000000000000000;
		num2 = 32'b00111111110000000000000000000000;
		func = 3'b011;
 //8.25/1.5=5.5 01000000101100000000000000000000
		
		#10;
		// div test 
      num1 = 32'b11000001000001000000000000000000;
		num2 = 32'b00111111110000000000000000000000;
		func = 3'b011;
 //-8.25/1.5=-5.5 11000000101100000000000000000000
 
		#10;
		// div over flow test 
      num1 = 32'b1_11111110_00001000000000000000000;
		num2 = 32'b0_00000001_10000000000000000000000;
		func = 3'b011;
 //over flow
		
	
		#10;
		// div inexact test 
      num1 = 32'b11000001000001000000000000000000;
		num2 = 32'b10111111101000000000000000000000;
		func = 3'b011;
 //-8.25/1.25=6.6 inexact 11000000101100000000000000000000
		
		
		#10;
		// div Qnan test 
      num1 = 32'b1_11111111_00000000000000000000000;
		num2 = 32'b0_11111111_00000000000000000000000;
		func = 3'b011;
 //Qnan
 
		#10;
		// inv test 
      num1 = 32'b01000000000000000000000000000000;
		num2 = 32'b0_11111111_00000000000000000000000;
		func = 3'b101;
 //1/2 = 0.5  00111111000000000000000000000000
 
		#10;
		// inv test 
      num1 = 32'b01000000000000000000000000000000;
		num2 = 32'b0_11111111_00000000000000000000000;
		func = 3'b101;
 //1/2 = 0.5  00111111000000000000000000000000
 
		#10;
		// inv div_by_zero test 
      num1 = 32'b00000000000000000000000000000000;
		num2 = 32'b0_11111111_00000000000000000000000;
		func = 3'b101;
 //1/0 = 0.5  div_by_zero
		
		#10;
		// div test 
      num1 = 32'b01111111100000000000000000000000;
		num2 = 32'b00111111110000000000000000000000;
		func = 3'b011;
 //inf/1.5=inf 01000000101100000000000000000000
 
		
		#10;
		// div test 
      num2 = 32'b01111111100000000000000000000000;
		num1 = 32'b00111111110000000000000000000000;
		func = 3'b011;
 //1.5/inf=0 01000000101100000000000000000000
		#10;
		// rounding test 
      num1 = 32'b01000000000000000000000000000000;
		num2 = 32'b0_11111111_00000000000000000000000;
		func = 3'b110;
 //2 = 2  01000000000000000000000000000000
 
		#10;
		// rounding test 
      num1 = 32'b01000000001000000000000000000000;
		num2 = 32'b0_11111111_00000000000000000000000;
		func = 3'b110;
 //2.5 = 3  01000000000000000000000000000000
		#10;
		// rounding test 
      num1 = 32'b11000000000100000000000000000000;
		num2 = 32'b0_11111111_00000000000000000000000;
		func = 3'b110;
 //-2.25 = -2  01000000000000000000000000000000
		#10
		// rounding overflow test 
      num1 = 32'b11111110000100000000000000000000;
		num2 = 32'b0_11111111_00000000000000000000000;
		func = 3'b110;
 //overflow  01000000000000000000000000000000
 
		
		#10;
		// rounding test 
      num1 = 32'b00111110100000000000000000000000;
		num2 = 32'b0_11111111_00000000000000000000000;
		func = 3'b110;
 //0.25 = 0  00000000000000000000000000000000
 
		#10;
		// cmp test 
      num1 = 32'b01000001000001000000000000000000;
		num2 = 32'b00111111110000000000000000000000;
		func = 3'b100;
 //8.25 > 1.5 = 001
		
		#10;
		// cmp test 
      num1 = 32'b11000001000001000000000000000000;
		num2 = 32'b00111111110000000000000000000000;
		func = 3'b100;
 //-8.25 < 1.5 = 100
		
		#10;
		// cmp test 
      num1 = 32'b11000001000001000000000000000000;
		num2 = 32'b10111111110000000000000000000000;
		func = 3'b100;
 //-8.25 < -1.5 = 100
		
		#10;
		// cmp test 
      num1 = 32'b11000001000001000000000000000000;
		num2 = 32'b11000001000001000000000000000000;
		func = 3'b100;
 //-8.25 == -8.25 = 010
		
		// Add stimulus here
  #10;    	
		
	end
       
endmodule

